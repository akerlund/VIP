////////////////////////////////////////////////////////////////////////////////
//
// Copyright (C) 2020 Fredrik Åkerlund
// https://github.com/akerlund/VIP
//
// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <https://www.gnu.org/licenses/>.
//
// Description:
//
////////////////////////////////////////////////////////////////////////////////

class clk_rst_config extends uvm_object;

  realtime clock_period      = 10.0;
  logic    rst_event_enabled = '0;

  `uvm_object_utils_begin(clk_rst_config);
  `uvm_field_real(clock_period,     UVM_DEFAULT)
  `uvm_field_int(rst_event_enabled, UVM_DEFAULT)
  `uvm_object_utils_end;

  function new(string name = "clk_rst_config");
    super.new(name);
  endfunction

endclass
