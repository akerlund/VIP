////////////////////////////////////////////////////////////////////////////////
//
// Copyright (C) 2021 Fredrik Åkerlund
//
// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <https://www.gnu.org/licenses/>.
//
// Description:
//
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
//                                                                            //
//           AUTOGENERATED FILE, DO NOT CHANGE THIS FILE MANUALLY.            //
//           CHANGE THE YAML FILE AND RERUN THE SCRIPT TO GENERATE.           //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////

// -----------------------------------------------------------------------------
// Command register
// -----------------------------------------------------------------------------
class command_reg extends uvm_reg;

  `uvm_object_utils(command_reg)

  rand uvm_reg_field cmd_command;


  function new (string name = "command_reg");
    super.new(name, 1, UVM_NO_COVERAGE);
  endfunction


  function void build();


    // -----------------------------------------------------------------------------
    // Command bit
    // -----------------------------------------------------------------------------
    cmd_command = uvm_reg_field::type_id::create("cmd_command");
    cmd_command.configure(
      .parent(this),
      .size(1),
      .lsb_pos(0),
      .access("WO"),
      .volatile(0),
      .reset(0),
      .has_reset(1),
      .is_rand(0),
      .individually_accessible(0)
    );
    add_hdl_path_slice("cmd_command", 0, 1);

  endfunction

endclass

// -----------------------------------------------------------------------------
// Configuration register
// -----------------------------------------------------------------------------
class configuration_reg extends uvm_reg;

  `uvm_object_utils(configuration_reg)

  rand uvm_reg_field cr_configuration;


  function new (string name = "configuration_reg");
    super.new(name, 64, UVM_NO_COVERAGE);
  endfunction


  function void build();


    // -----------------------------------------------------------------------------
    // Configuration register
    // -----------------------------------------------------------------------------
    cr_configuration = uvm_reg_field::type_id::create("cr_configuration");
    cr_configuration.configure(
      .parent(this),
      .size(64),
      .lsb_pos(0),
      .access("RW"),
      .volatile(0),
      .reset(0),
      .has_reset(1),
      .is_rand(0),
      .individually_accessible(0)
    );
    add_hdl_path_slice("cr_configuration", 0, 64);

  endfunction

endclass

// -----------------------------------------------------------------------------
// Status register
// -----------------------------------------------------------------------------
class status_reg extends uvm_reg;

  `uvm_object_utils(status_reg)

  rand uvm_reg_field sr_status;


  function new (string name = "status_reg");
    super.new(name, 64, UVM_NO_COVERAGE);
  endfunction


  function void build();


    // -----------------------------------------------------------------------------
    // Status register
    // -----------------------------------------------------------------------------
    sr_status = uvm_reg_field::type_id::create("sr_status");
    sr_status.configure(
      .parent(this),
      .size(64),
      .lsb_pos(0),
      .access("RW"),
      .volatile(0),
      .reset(0),
      .has_reset(0),
      .is_rand(0),
      .individually_accessible(0)
    );
    add_hdl_path_slice("sr_status", 0, 64);

  endfunction

endclass

