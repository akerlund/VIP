////////////////////////////////////////////////////////////////////////////////
//
// Copyright (C) 2021 Fredrik Åkerlund
// https://github.com/akerlund/VIP
//
// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <https://www.gnu.org/licenses/>.
//
// Description:
//
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
//                                                                            //
//           AUTOGENERATED FILE, DO NOT CHANGE THIS FILE MANUALLY.            //
//           CHANGE THE YAML FILE AND RERUN THE SCRIPT TO GENERATE.           //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////


import axi4_address_pkg::*;

module axi4_axi_slave #(
    parameter int AXI_ADDR_WIDTH_P = -1,
    parameter int AXI_DATA_WIDTH_P = -1,
    parameter int AXI_ID_P = -1
  )(
    axi_cfg_if.slave cif,
    output logic          cmd_command,
    output logic [63 : 0] cr_configuration,
    input  wire  [63 : 0] sr_status
  );

  localparam logic [1 : 0] AXI_RESP_SLVERR_C = 2'b01;

  // ---------------------------------------------------------------------------
  // Internal signals
  // ---------------------------------------------------------------------------

  typedef enum {
    WAIT_MST_AWVALID_E,
    WAIT_FOR_BREADY_E,
    WAIT_MST_WLAST_E
  } write_state_t;

  write_state_t write_state;

  logic [AXI_ADDR_WIDTH_P-1 : 0] awaddr_r0;

  typedef enum {
    WAIT_MST_ARVALID_E,
    WAIT_SLV_RLAST_E
  } read_state_t;

  read_state_t read_state;

  logic [AXI_ADDR_WIDTH_P-1 : 0] araddr_r0;
  logic                  [7 : 0] arlen_c0;
  logic                  [7 : 0] arlen_r0;
  logic [AXI_DATA_WIDTH_P-1 : 0] rdata_c0;
  logic                  [1 : 0] rresp_c0;



  // ---------------------------------------------------------------------------
  // Port assignments
  // ---------------------------------------------------------------------------

  assign cif.rid = AXI_ID_P;

  // ---------------------------------------------------------------------------
  // Write processes
  // ---------------------------------------------------------------------------
  always_ff @(posedge cif.clk or negedge cif.rst_n) begin
    if (!cif.rst_n) begin

      write_state <= WAIT_MST_AWVALID_E;
      awaddr_r0   <= '0;
      cif.awready <= '0;
      cif.wready  <= '0;
      cif.bid     <= '0;
      cif.bvalid  <= '0;
      cif.bresp   <= '0;
      cmd_command      <= 0;
      cr_configuration <= 0;

    end
    else begin

      cmd_command <= '0;



      case (write_state)

        default: begin
          write_state <= WAIT_MST_AWVALID_E;
        end

        WAIT_MST_AWVALID_E: begin

          cif.awready <= '1;

          if (cif.awvalid && cif.awready) begin
            write_state <= WAIT_MST_WLAST_E;
            cif.awready <= '0;
            cif.bid     <= cif.awid;
            awaddr_r0   <= cif.awaddr;
            cif.wready  <= '1;
          end

        end


        WAIT_FOR_BREADY_E: begin

          if (cif.bvalid && cif.bready) begin
            write_state <= WAIT_MST_AWVALID_E;
            cif.awready <= '1;
            cif.bvalid  <= '0;
            cif.bresp   <= '0;
          end

        end


        WAIT_MST_WLAST_E: begin

          if (cif.wlast && cif.wvalid) begin
            write_state <= WAIT_FOR_BREADY_E;
            cif.bvalid  <= '1;
            cif.wready  <= '0;
          end


          if (cif.wvalid) begin

            awaddr_r0 <= awaddr_r0 + (AXI_DATA_WIDTH_P/8);

            case (awaddr_r0)

              COMMAND_ADDR: begin
                cmd_command <= cif.wdata[0];
              end

              CONFIGURATION_ADDR: begin
                cr_configuration <= cif.wdata[63 : 0];
              end


              default: begin
                cif.bresp <= AXI_RESP_SLVERR_C;
              end

            endcase


          end
        end
      endcase
    end
  end

  // ---------------------------------------------------------------------------
  // Read process
  // ---------------------------------------------------------------------------

  assign cif.rlast = cif.rvalid && arlen_r0 == '0;

  always_comb begin
    arlen_c0 = arlen_r0;

    case (read_state)
      WAIT_MST_ARVALID_E: begin
        if (cif.arvalid && cif.arready) begin
          arlen_c0 = cif.arlen;
        end
      end

      WAIT_SLV_RLAST_E: begin
        if (cif.rready && cif.rvalid) begin
          if (arlen_r0 != '0) begin
            arlen_c0 = arlen_r0 - 1;
          end
        end
      end
    endcase
  end

  // FSM
  always_ff @(posedge cif.clk or negedge cif.rst_n) begin
    if (!cif.rst_n) begin

      read_state  <= WAIT_MST_ARVALID_E;
      cif.arready <= '0;
      araddr_r0   <= '0;
      arlen_r0    <= '0;
      cif.rid     <= '0;
      cif.rdata   <= '0;
      cif.rresp   <= '0;
      cif.rvalid  <= '0;

    end
    else begin

      case (read_state)

        default: begin
          read_state <= WAIT_MST_ARVALID_E;
        end

        WAIT_MST_ARVALID_E: begin

          cif.arready <= '1;

          if (cif.arvalid && cif.arready) begin
            read_state  <= WAIT_SLV_RLAST_E;
            araddr_r0   <= cif.araddr;
            cif.rid     <= cif.arid;
            cif.arready <= '0;
          end

        end

        WAIT_SLV_RLAST_E: begin

          cif.rvalid <= '1;
          cif.rdata  <= rdata_c0;
          cif.rresp  <= rresp_c0;

          if (cif.rready && cif.rvalid) begin
            araddr_r0 <= araddr_r0 + (AXI_DATA_WIDTH_P/8);
          end

          if (cif.rvalid && cif.rready && cif.rlast) begin
            read_state  <= WAIT_MST_ARVALID_E;
            cif.arready <= '1;
            cif.rvalid  <= '0;
          end

        end
      endcase
    end
  end



  always_comb begin

    rdata_c0 = '0;
    rresp_c0 = '0;

    case (araddr_r0)

      CONFIGURATION_ADDR: begin
        rdata_c0 = cr_configuration;
      end

      STATUS_ADDR: begin
        rdata_c0 = sr_status;
      end

      default: begin
        rresp_c0 = AXI_RESP_SLVERR_C;
        rdata_c0 = '0;
      end

    endcase
  end

endmodule
