////////////////////////////////////////////////////////////////////////////////
//
// Copyright (C) 2021 Fredrik Åkerlund
// https://github.com/akerlund/VIP
//
// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <https://www.gnu.org/licenses/>.
//
// Description:
//
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
//                                                                            //
//           AUTOGENERATED FILE, DO NOT CHANGE THIS FILE MANUALLY.            //
//           CHANGE THE YAML FILE AND RERUN THE SCRIPT TO GENERATE.           //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////


`ifndef AXI4_ADDRESS_PKG
`define AXI4_ADDRESS_PKG

package axi4_address_pkg;

  localparam logic [15 : 0] AXI4_HIGH_ADDRESS  = 16'h0018;
  localparam logic [15 : 0] COMMAND_ADDR       = 16'h0000;
  localparam logic [15 : 0] CONFIGURATION_ADDR = 16'h0008;
  localparam logic [15 : 0] STATUS_ADDR        = 16'h0010;

endpackage

`endif
