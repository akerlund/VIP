////////////////////////////////////////////////////////////////////////////////
//
// Copyright (C) 2021 Fredrik Åkerlund
// https://github.com/akerlund/VIP
//
// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <https://www.gnu.org/licenses/>.
//
// Description:
//
////////////////////////////////////////////////////////////////////////////////

class vip_axi4_monitor_callback extends uvm_callback;

  `uvm_object_utils(vip_axi4_monitor_callback)

  function new(string name = "vip_axi4_monitor_callback");
    super.new(name);
  endfunction

  task pre_drive;
    //`uvm_info("USER_CALLBACK","Inside pre_drive method",UVM_LOW);
  endtask
  task post_drive;
    //`uvm_info("USER_CALLBACK","Inside post_drive method",UVM_LOW);
  endtask

  endclass
